netcdf domain_input {
dimensions:
        x = 5 ;
        y = 5 ;
        x_resample = 2 ;
        y_resample = 2 ;
	nbounds = 2 ;
variables:
        float x(x) ;
                x:long_name = "original x coordinate" ;
                x:units = "1";
		x:bounds = "x_bounds" ;
        float y(y) ;
                y:long_name = "original y coordinate" ;
                y:units = "1";
                y:bounds = "y_bounds" ;
        float x_resample(x_resample) ;
                x_resample:long_name = "resampled x coordinate" ;
                x_resample:units = "1";
		x_resample:bounds = "x_resample_bounds" ;
        float y_resample(y_resample) ;
                y_resample:long_name = "resampled y coordinate" ;
                y_resample:units = "1";
		y_resample:bounds = "y_resample_bounds";
	float x_bounds(x, nbounds) ;
	float y_bounds(y, nbounds) ;
	float x_resample_bounds(x_resample, nbounds) ;
	float y_resample_bounds(y_resample, nbounds) ;
        double original_data(y,x) ;
                original_data:long_name = "input data values" ;
                original_data:units = "1";
        double resample_data(y_resample,x_resample) ;
                resample_data:long_name = "expected resampled data values" ;
                resample_data:units = "1";

// global attributes:
                :title = "Input data for XIOS Domain resampling; data is a sum of the x & y coordinates; x + y ." ;

data:

 x = 0, 2, 4, 6, 8 ;

 y = 0, 2, 4, 6, 8 ;

 x_resample = 3, 5 ;

 y_resample = 3, 5 ;

 x_bounds = -1, 1, 1, 3, 3, 5, 5, 7, 7, 9 ;

 y_bounds = -1, 1, 1, 3, 3, 5, 5, 7, 7, 9 ;

 x_resample_bounds = 2, 4, 4, 6 ;

 y_resample_bounds = 2, 4, 4, 6 ;

 original_data =  0,  2,  4,  6,  8,
                  2,  4,  6,  8, 10,
                  4,  6,  8, 10, 12,
                  6,  8, 10, 12, 14,
                  8, 10, 12, 14, 16 ;

 resample_data = 6, 8,
                 8, 10 ;

}
